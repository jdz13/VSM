@Filename: C:\vsm-lv\Jake\Angles\Minor loops\SP6772\SP6772_minor-a000-00.VHD
@Measurement Controlfilename: C:\vsm-lv\Reinoud\Recipes\Jake\Angles\SP6772_minor-a000-00.VHC
@Calibration filename: c:\vsm-lv\Reinoud\settings\default.cal
@Parameter Filec:\vsm-lv\Reinoud\settings\default.cal
@Operator: Reinoud
@Samplename: SP6772
@Date: Wednesday, July 18, 2018    (2018-07-18)
@Time: 15:52:50
@Test ID: test
@Apparatus: EV X; SN: XXXXXXXX; Customer: XXXXXXXXX; first started on: Tuesday, January 25, 2011
VSM Model = EV X, Signal Processor = 2 SRS SR 830, Gaussmeter = 32 KP DRC, Gauss Probe = 1 x, VSM = TRUE, Torque = FALSE
Rotation Card = TRUE, Rotation Display = FALSE, Rotate Option = Mdrive
Temperature Control = TRUE, Temperature control Type = SI 9700, Thermocouple Type = J-type, Liquid Helium = FALSE, Boil Off Nitrogen = FALSE, Leave Temp On = FALSE
Vector Coils = TRUE, Z Coils = FALSE, Stationary Coils = FALSE, Sensor Angle = 0 deg, Signal Connection = A-B
@System Status = Online
@Sample Orientation and Shape: line parallel with field
@@Sample Dimensions
Shape = Circular;  Length = 6.60 [mm] Width = 6.60 [mm] Thickness = 1.000E+3 [nm] Diameter = 8.00 [mm] Volume : 5.027E-11 [m^3] Area = 5.027E+1 [mm^2] Mass = 1.000E+0 [g] Nd =  0.00 Sample Angle Offset = 0.000 
Ms (for Hys loss calculation) = 1.000 [memu]
@@End Sample Dimensions
@Measurement type: Hysteresis Loop
@Product of: MicroSense EasyVSM Software version 9.13U (January 27, 2011)
@@Comments: 
@@END Comments
@@Parameters
@@Measurement Preparation Actions
Action 0:      Set Field Angle to 0.0000 [deg] and wait 0.0000 s ; Set Mode = Set and wait till there
@@END Measurement Preparation Actions
@@Measurement Parameters
@Repeat all sections = Symmetric
@Number of sections= 7
@Section 0: Hysteresis; New Plot
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Repeated Actions:
Action 0:      Set Applied Field to 0.0000 [Oe] and wait 0.0000 s ; Set Mode = Set and wait till there; Measure 
@Main Parameter = 0 : Applied Field [Oe].
@Main Parameter Setup:
     From: -17000.0000 [Oe] To: -1000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Measured Signal(s) = X
@Section 0 END
@Section 1: Hysteresis
@Preparation Actions:
Action 0:      Set Gauss Range to 1.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Main Parameter Setup:
     From: -1000.0000 [Oe] To: -500.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 1 END
@Section 2: Hysteresis
@Main Parameter Setup:
     From: -500.0000 [Oe] To: -100.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 2 END
@Section 3: Hysteresis
@Preparation Actions:
Action 0:      Set Gauss Range to 2.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Main Parameter Setup:
     From: -100.0000 [Oe] To: 100.0000 [Oe] Min Stepsize/Sweeprate = 10.0000 [Oe] Max Stepsize/Sweeprate = 10.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 3 END
@Section 4: Hysteresis
@Preparation Actions:
Action 0:      Set Gauss Range to 1.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Main Parameter Setup:
     From: 100.0000 [Oe] To: 500.0000 [Oe] Min Stepsize/Sweeprate = 50.0000 [Oe] Max Stepsize/Sweeprate = 50.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 4 END
@Section 5: Hysteresis
@Main Parameter Setup:
     From: 500.0000 [Oe] To: 1000.0000 [Oe] Min Stepsize/Sweeprate = 100.0000 [Oe] Max Stepsize/Sweeprate = 100.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 5 END
@Section 6: Hysteresis
@Preparation Actions:
Action 0:      Set Gauss Range to 0.0000 [ ] and wait 0.0000 s ; Set Mode = Set and wait till there
@Main Parameter Setup:
     From: 1000.0000 [Oe] To: 17000.0000 [Oe] Min Stepsize/Sweeprate = 1000.0000 [Oe] Max Stepsize/Sweeprate = 1000.0000 [Oe]
     Signal change min step =  0.00 [%] Signal change max step =  0.00 [%] ;  Wait time =    0.00 [sec] Up & Down = No
@Section 6 END
@@Plot Settings
Number of plots: 1
Plot 0: Hysteresis = On; Section: 0; Signal: X; Label: Hys X; Point style: 1; Interpolation: On; Color: 16777222; Mirror: Off
@@ENDPlot Settings
@@END Measurement Parameters
@@Instrument Parameters
Stationary Coils = FALSE
Sensor Angle = 0 deg
@Gauss Range: 30 kOe
@Emu Range: 1 mV
@Torque Range: 4000 dyne cm
@Auto-range emu: No
@Number of averages: 10
@Rot 0 deg cal: -21000
@Rot 360 deg cal: 21000
@Dec Pt. constant: 1000
@Emu dec cal: 100
@Emdac: 28000
@Emu/v: 72.879
@Y Coils Correction Factor: 1.440
@Sample Shape Correction Factor: 1.000
@Coil Angle Alpha: 45.000
@Coil Angle Beta: -45.000
[Data Manipulation]
Field Linearity Correction = No
Image Effect Correction = Yes
Image Correction Array Length = 21
12499.000000   1.000000
12748.000000   0.999735
12998.000000   0.999575
13249.000000   0.999364
13499.000000   0.999258
13749.000000   0.999205
13999.000000   0.999100
14248.000000   0.999100
14498.000000   0.999205
14748.000000   0.999312
14998.000000   0.999417
15248.000000   0.999682
15499.000000   0.999840
15748.000000   1.000106
15999.000000   1.000424
16248.000000   1.000795
16498.000000   1.001166
16748.000000   1.001697
16998.000000   1.002176
17248.000000   1.002708
17498.000000   1.003401
Sample image effect correction factor = 1.000000, Sample holder image effect correction factor = 1.000000
Background Subtraction = Yes   Method = Straight Line
Background slope x, y, z [emu/Oe] = -6.188366E-8   -2.604465E-9   0.000000E+0
Background Offset x, y, z [emu] = -9.024043E-6   5.450853E-6   0.000000E+0
Angular Sensitivity Correction = Yes
Angular Sensitivity array length = 361
0.000000   9.995411E-1   1.478461E+0   0.000000
1.000000   9.974509E-1   1.478734E+0   0.000000
2.000000   9.953678E-1   1.479006E+0   0.000000
3.000000   9.932991E-1   1.479275E+0   0.000000
4.000000   9.912518E-1   1.479539E+0   0.000000
5.000000   9.892331E-1   1.479797E+0   0.000000
6.000000   9.872502E-1   1.480047E+0   0.000000
7.000000   9.853102E-1   1.480288E+0   0.000000
8.000000   9.834203E-1   1.480518E+0   0.000000
9.000000   9.815877E-1   1.480735E+0   0.000000
10.000000   9.798194E-1   1.480939E+0   0.000000
11.000000   9.781226E-1   1.481127E+0   0.000000
12.000000   9.765046E-1   1.481298E+0   0.000000
13.000000   9.749724E-1   1.481450E+0   0.000000
14.000000   9.735332E-1   1.481582E+0   0.000000
15.000000   9.721941E-1   1.481692E+0   0.000000
16.000000   9.709610E-1   1.481777E+0   0.000000
17.000000   9.698342E-1   1.481826E+0   0.000000
18.000000   9.688126E-1   1.481825E+0   0.000000
19.000000   9.678951E-1   1.481761E+0   0.000000
20.000000   9.670809E-1   1.481622E+0   0.000000
21.000000   9.663687E-1   1.481393E+0   0.000000
22.000000   9.657576E-1   1.481063E+0   0.000000
23.000000   9.652465E-1   1.480617E+0   0.000000
24.000000   9.648345E-1   1.480042E+0   0.000000
25.000000   9.645203E-1   1.479326E+0   0.000000
26.000000   9.643031E-1   1.478456E+0   0.000000
27.000000   9.641818E-1   1.477417E+0   0.000000
28.000000   9.641553E-1   1.476198E+0   0.000000
29.000000   9.642226E-1   1.474784E+0   0.000000
30.000000   9.643826E-1   1.473164E+0   0.000000
31.000000   9.646346E-1   1.471326E+0   0.000000
32.000000   9.649784E-1   1.469273E+0   0.000000
33.000000   9.654142E-1   1.467010E+0   0.000000
34.000000   9.659421E-1   1.464542E+0   0.000000
35.000000   9.665623E-1   1.461875E+0   0.000000
36.000000   9.672748E-1   1.459015E+0   0.000000
37.000000   9.680799E-1   1.455965E+0   0.000000
38.000000   9.689777E-1   1.452732E+0   0.000000
39.000000   9.699683E-1   1.449320E+0   0.000000
40.000000   9.710519E-1   1.445736E+0   0.000000
41.000000   9.722285E-1   1.441983E+0   0.000000
42.000000   9.734984E-1   1.438069E+0   0.000000
43.000000   9.748616E-1   1.433997E+0   0.000000
44.000000   9.763183E-1   1.429773E+0   0.000000
45.000000   9.778686E-1   1.425402E+0   0.000000
46.000000   9.795120E-1   1.420891E+0   0.000000
47.000000   9.812448E-1   1.416248E+0   0.000000
48.000000   9.830627E-1   1.411485E+0   0.000000
49.000000   9.849614E-1   1.406611E+0   0.000000
50.000000   9.869365E-1   1.401636E+0   0.000000
51.000000   9.889837E-1   1.396571E+0   0.000000
52.000000   9.910986E-1   1.391426E+0   0.000000
53.000000   9.932770E-1   1.386211E+0   0.000000
54.000000   9.955145E-1   1.380936E+0   0.000000
55.000000   9.978067E-1   1.375612E+0   0.000000
56.000000   1.000149E+0   1.370249E+0   0.000000
57.000000   1.002538E+0   1.364857E+0   0.000000
58.000000   1.004969E+0   1.359446E+0   0.000000
59.000000   1.007437E+0   1.354026E+0   0.000000
60.000000   1.009938E+0   1.348609E+0   0.000000
61.000000   1.012470E+0   1.343204E+0   0.000000
62.000000   1.015040E+0   1.337826E+0   0.000000
63.000000   1.017658E+0   1.332491E+0   0.000000
64.000000   1.020332E+0   1.327213E+0   0.000000
65.000000   1.023073E+0   1.322007E+0   0.000000
66.000000   1.025889E+0   1.316890E+0   0.000000
67.000000   1.028791E+0   1.311875E+0   0.000000
68.000000   1.031787E+0   1.306979E+0   0.000000
69.000000   1.034887E+0   1.302215E+0   0.000000
70.000000   1.038100E+0   1.297601E+0   0.000000
71.000000   1.041435E+0   1.293150E+0   0.000000
72.000000   1.044902E+0   1.288878E+0   0.000000
73.000000   1.048511E+0   1.284799E+0   0.000000
74.000000   1.052271E+0   1.280930E+0   0.000000
75.000000   1.056190E+0   1.277286E+0   0.000000
76.000000   1.060275E+0   1.273874E+0   0.000000
77.000000   1.064511E+0   1.270678E+0   0.000000
78.000000   1.068882E+0   1.267675E+0   0.000000
79.000000   1.073371E+0   1.264841E+0   0.000000
80.000000   1.077959E+0   1.262152E+0   0.000000
81.000000   1.082630E+0   1.259585E+0   0.000000
82.000000   1.087366E+0   1.257116E+0   0.000000
83.000000   1.092150E+0   1.254722E+0   0.000000
84.000000   1.096965E+0   1.252380E+0   0.000000
85.000000   1.101792E+0   1.250065E+0   0.000000
86.000000   1.106615E+0   1.247755E+0   0.000000
87.000000   1.111417E+0   1.245425E+0   0.000000
88.000000   1.116179E+0   1.243053E+0   0.000000
89.000000   1.120885E+0   1.240614E+0   0.000000
90.000000   1.125517E+0   1.238086E+0   0.000000
91.000000   1.130059E+0   1.235451E+0   0.000000
92.000000   1.134507E+0   1.232719E+0   0.000000
93.000000   1.138856E+0   1.229906E+0   0.000000
94.000000   1.143101E+0   1.227029E+0   0.000000
95.000000   1.147240E+0   1.224104E+0   0.000000
96.000000   1.151268E+0   1.221147E+0   0.000000
97.000000   1.155181E+0   1.218174E+0   0.000000
98.000000   1.158976E+0   1.215203E+0   0.000000
99.000000   1.162648E+0   1.212249E+0   0.000000
100.000000   1.166194E+0   1.209329E+0   0.000000
101.000000   1.169609E+0   1.206459E+0   0.000000
102.000000   1.172890E+0   1.203655E+0   0.000000
103.000000   1.176033E+0   1.200933E+0   0.000000
104.000000   1.179033E+0   1.198311E+0   0.000000
105.000000   1.181888E+0   1.195803E+0   0.000000
106.000000   1.184594E+0   1.193425E+0   0.000000
107.000000   1.187151E+0   1.191176E+0   0.000000
108.000000   1.189560E+0   1.189057E+0   0.000000
109.000000   1.191822E+0   1.187066E+0   0.000000
110.000000   1.193939E+0   1.185202E+0   0.000000
111.000000   1.195912E+0   1.183464E+0   0.000000
112.000000   1.197741E+0   1.181850E+0   0.000000
113.000000   1.199428E+0   1.180359E+0   0.000000
114.000000   1.200974E+0   1.178991E+0   0.000000
115.000000   1.202380E+0   1.177744E+0   0.000000
116.000000   1.203648E+0   1.176616E+0   0.000000
117.000000   1.204777E+0   1.175607E+0   0.000000
118.000000   1.205770E+0   1.174715E+0   0.000000
119.000000   1.206627E+0   1.173940E+0   0.000000
120.000000   1.207349E+0   1.173280E+0   0.000000
121.000000   1.207939E+0   1.172734E+0   0.000000
122.000000   1.208399E+0   1.172305E+0   0.000000
123.000000   1.208732E+0   1.171996E+0   0.000000
124.000000   1.208942E+0   1.171809E+0   0.000000
125.000000   1.209032E+0   1.171747E+0   0.000000
126.000000   1.209007E+0   1.171813E+0   0.000000
127.000000   1.208868E+0   1.172009E+0   0.000000
128.000000   1.208620E+0   1.172339E+0   0.000000
129.000000   1.208266E+0   1.172805E+0   0.000000
130.000000   1.207809E+0   1.173411E+0   0.000000
131.000000   1.207253E+0   1.174158E+0   0.000000
132.000000   1.206602E+0   1.175050E+0   0.000000
133.000000   1.205858E+0   1.176090E+0   0.000000
134.000000   1.205025E+0   1.177279E+0   0.000000
135.000000   1.204107E+0   1.178622E+0   0.000000
136.000000   1.203105E+0   1.180119E+0   0.000000
137.000000   1.202012E+0   1.181762E+0   0.000000
138.000000   1.200819E+0   1.183543E+0   0.000000
139.000000   1.199519E+0   1.185452E+0   0.000000
140.000000   1.198102E+0   1.187481E+0   0.000000
141.000000   1.196559E+0   1.189620E+0   0.000000
142.000000   1.194883E+0   1.191859E+0   0.000000
143.000000   1.193063E+0   1.194190E+0   0.000000
144.000000   1.191092E+0   1.196604E+0   0.000000
145.000000   1.188961E+0   1.199092E+0   0.000000
146.000000   1.186661E+0   1.201643E+0   0.000000
147.000000   1.184184E+0   1.204250E+0   0.000000
148.000000   1.181520E+0   1.206902E+0   0.000000
149.000000   1.178662E+0   1.209592E+0   0.000000
150.000000   1.175600E+0   1.212309E+0   0.000000
151.000000   1.172327E+0   1.215048E+0   0.000000
152.000000   1.168848E+0   1.217818E+0   0.000000
153.000000   1.165167E+0   1.220632E+0   0.000000
154.000000   1.161288E+0   1.223503E+0   0.000000
155.000000   1.157217E+0   1.226442E+0   0.000000
156.000000   1.152959E+0   1.229464E+0   0.000000
157.000000   1.148519E+0   1.232580E+0   0.000000
158.000000   1.143902E+0   1.235803E+0   0.000000
159.000000   1.139113E+0   1.239147E+0   0.000000
160.000000   1.134157E+0   1.242622E+0   0.000000
161.000000   1.129038E+0   1.246243E+0   0.000000
162.000000   1.123763E+0   1.250022E+0   0.000000
163.000000   1.118335E+0   1.253972E+0   0.000000
164.000000   1.112761E+0   1.258104E+0   0.000000
165.000000   1.107045E+0   1.262433E+0   0.000000
166.000000   1.101194E+0   1.266966E+0   0.000000
167.000000   1.095231E+0   1.271691E+0   0.000000
168.000000   1.089177E+0   1.276593E+0   0.000000
169.000000   1.083057E+0   1.281656E+0   0.000000
170.000000   1.076894E+0   1.286865E+0   0.000000
171.000000   1.070713E+0   1.292202E+0   0.000000
172.000000   1.064535E+0   1.297653E+0   0.000000
173.000000   1.058386E+0   1.303202E+0   0.000000
174.000000   1.052288E+0   1.308833E+0   0.000000
175.000000   1.046265E+0   1.314529E+0   0.000000
176.000000   1.040340E+0   1.320275E+0   0.000000
177.000000   1.034538E+0   1.326056E+0   0.000000
178.000000   1.028881E+0   1.331855E+0   0.000000
179.000000   1.023394E+0   1.337656E+0   0.000000
180.000000   1.018099E+0   1.343444E+0   0.000000
181.000000   1.013016E+0   1.349202E+0   0.000000
182.000000   1.008143E+0   1.354916E+0   0.000000
183.000000   1.003473E+0   1.360569E+0   0.000000
184.000000   9.990010E-1   1.366147E+0   0.000000
185.000000   9.947191E-1   1.371632E+0   0.000000
186.000000   9.906216E-1   1.377011E+0   0.000000
187.000000   9.867020E-1   1.382266E+0   0.000000
188.000000   9.829538E-1   1.387384E+0   0.000000
189.000000   9.793706E-1   1.392347E+0   0.000000
190.000000   9.759461E-1   1.397140E+0   0.000000
191.000000   9.726738E-1   1.401749E+0   0.000000
192.000000   9.695473E-1   1.406157E+0   0.000000
193.000000   9.665602E-1   1.410348E+0   0.000000
194.000000   9.637061E-1   1.414307E+0   0.000000
195.000000   9.609785E-1   1.418019E+0   0.000000
196.000000   9.583727E-1   1.421472E+0   0.000000
197.000000   9.558905E-1   1.424669E+0   0.000000
198.000000   9.535352E-1   1.427616E+0   0.000000
199.000000   9.513104E-1   1.430322E+0   0.000000
200.000000   9.492193E-1   1.432794E+0   0.000000
201.000000   9.472655E-1   1.435038E+0   0.000000
202.000000   9.454524E-1   1.437061E+0   0.000000
203.000000   9.437833E-1   1.438871E+0   0.000000
204.000000   9.422618E-1   1.440476E+0   0.000000
205.000000   9.408912E-1   1.441881E+0   0.000000
206.000000   9.396749E-1   1.443094E+0   0.000000
207.000000   9.386164E-1   1.444122E+0   0.000000
208.000000   9.377190E-1   1.444973E+0   0.000000
209.000000   9.369863E-1   1.445653E+0   0.000000
210.000000   9.364216E-1   1.446170E+0   0.000000
211.000000   9.360260E-1   1.446530E+0   0.000000
212.000000   9.357914E-1   1.446744E+0   0.000000
213.000000   9.357072E-1   1.446820E+0   0.000000
214.000000   9.357631E-1   1.446766E+0   0.000000
215.000000   9.359484E-1   1.446594E+0   0.000000
216.000000   9.362528E-1   1.446310E+0   0.000000
217.000000   9.366656E-1   1.445926E+0   0.000000
218.000000   9.371766E-1   1.445449E+0   0.000000
219.000000   9.377751E-1   1.444889E+0   0.000000
220.000000   9.384506E-1   1.444256E+0   0.000000
221.000000   9.391928E-1   1.443558E+0   0.000000
222.000000   9.399911E-1   1.442804E+0   0.000000
223.000000   9.408350E-1   1.442005E+0   0.000000
224.000000   9.417140E-1   1.441168E+0   0.000000
225.000000   9.426177E-1   1.440303E+0   0.000000
226.000000   9.435393E-1   1.439415E+0   0.000000
227.000000   9.444873E-1   1.438494E+0   0.000000
228.000000   9.454738E-1   1.437523E+0   0.000000
229.000000   9.465110E-1   1.436488E+0   0.000000
230.000000   9.476111E-1   1.435374E+0   0.000000
231.000000   9.487862E-1   1.434165E+0   0.000000
232.000000   9.500486E-1   1.432847E+0   0.000000
233.000000   9.514103E-1   1.431405E+0   0.000000
234.000000   9.528837E-1   1.429822E+0   0.000000
235.000000   9.544808E-1   1.428084E+0   0.000000
236.000000   9.562138E-1   1.426177E+0   0.000000
237.000000   9.580950E-1   1.424084E+0   0.000000
238.000000   9.601365E-1   1.421791E+0   0.000000
239.000000   9.623504E-1   1.419282E+0   0.000000
240.000000   9.647490E-1   1.416543E+0   0.000000
241.000000   9.673407E-1   1.413562E+0   0.000000
242.000000   9.701195E-1   1.410344E+0   0.000000
243.000000   9.730753E-1   1.406899E+0   0.000000
244.000000   9.761985E-1   1.403236E+0   0.000000
245.000000   9.794791E-1   1.399363E+0   0.000000
246.000000   9.829073E-1   1.395291E+0   0.000000
247.000000   9.864733E-1   1.391028E+0   0.000000
248.000000   9.901672E-1   1.386582E+0   0.000000
249.000000   9.939791E-1   1.381965E+0   0.000000
250.000000   9.978993E-1   1.377184E+0   0.000000
251.000000   1.001918E+0   1.372248E+0   0.000000
252.000000   1.006025E+0   1.367168E+0   0.000000
253.000000   1.010211E+0   1.361951E+0   0.000000
254.000000   1.014465E+0   1.356608E+0   0.000000
255.000000   1.018779E+0   1.351147E+0   0.000000
256.000000   1.023140E+0   1.345580E+0   0.000000
257.000000   1.027530E+0   1.339933E+0   0.000000
258.000000   1.031928E+0   1.334232E+0   0.000000
259.000000   1.036314E+0   1.328504E+0   0.000000
260.000000   1.040668E+0   1.322779E+0   0.000000
261.000000   1.044968E+0   1.317082E+0   0.000000
262.000000   1.049195E+0   1.311442E+0   0.000000
263.000000   1.053329E+0   1.305886E+0   0.000000
264.000000   1.057348E+0   1.300441E+0   0.000000
265.000000   1.061233E+0   1.295136E+0   0.000000
266.000000   1.064963E+0   1.289997E+0   0.000000
267.000000   1.068517E+0   1.285052E+0   0.000000
268.000000   1.071876E+0   1.280328E+0   0.000000
269.000000   1.075018E+0   1.275854E+0   0.000000
270.000000   1.077924E+0   1.271656E+0   0.000000
271.000000   1.080579E+0   1.267756E+0   0.000000
272.000000   1.082996E+0   1.264149E+0   0.000000
273.000000   1.085193E+0   1.260823E+0   0.000000
274.000000   1.087190E+0   1.257766E+0   0.000000
275.000000   1.089004E+0   1.254967E+0   0.000000
276.000000   1.090656E+0   1.252414E+0   0.000000
277.000000   1.092164E+0   1.250097E+0   0.000000
278.000000   1.093546E+0   1.248003E+0   0.000000
279.000000   1.094821E+0   1.246121E+0   0.000000
280.000000   1.096008E+0   1.244439E+0   0.000000
281.000000   1.097127E+0   1.242946E+0   0.000000
282.000000   1.098195E+0   1.241630E+0   0.000000
283.000000   1.099231E+0   1.240480E+0   0.000000
284.000000   1.100255E+0   1.239484E+0   0.000000
285.000000   1.101285E+0   1.238631E+0   0.000000
286.000000   1.102336E+0   1.237911E+0   0.000000
287.000000   1.103401E+0   1.237323E+0   0.000000
288.000000   1.104471E+0   1.236867E+0   0.000000
289.000000   1.105536E+0   1.236544E+0   0.000000
290.000000   1.106587E+0   1.236355E+0   0.000000
291.000000   1.107612E+0   1.236300E+0   0.000000
292.000000   1.108603E+0   1.236379E+0   0.000000
293.000000   1.109549E+0   1.236594E+0   0.000000
294.000000   1.110440E+0   1.236945E+0   0.000000
295.000000   1.111267E+0   1.237433E+0   0.000000
296.000000   1.112019E+0   1.238058E+0   0.000000
297.000000   1.112687E+0   1.238821E+0   0.000000
298.000000   1.113260E+0   1.239722E+0   0.000000
299.000000   1.113729E+0   1.240762E+0   0.000000
300.000000   1.114084E+0   1.241941E+0   0.000000
301.000000   1.114315E+0   1.243260E+0   0.000000
302.000000   1.114420E+0   1.244710E+0   0.000000
303.000000   1.114395E+0   1.246284E+0   0.000000
304.000000   1.114237E+0   1.247972E+0   0.000000
305.000000   1.113945E+0   1.249768E+0   0.000000
306.000000   1.113516E+0   1.251661E+0   0.000000
307.000000   1.112947E+0   1.253645E+0   0.000000
308.000000   1.112235E+0   1.255710E+0   0.000000
309.000000   1.111378E+0   1.257848E+0   0.000000
310.000000   1.110372E+0   1.260051E+0   0.000000
311.000000   1.109217E+0   1.262310E+0   0.000000
312.000000   1.107908E+0   1.264617E+0   0.000000
313.000000   1.106444E+0   1.266964E+0   0.000000
314.000000   1.104821E+0   1.269341E+0   0.000000
315.000000   1.103038E+0   1.271742E+0   0.000000
316.000000   1.101093E+0   1.274160E+0   0.000000
317.000000   1.098996E+0   1.276610E+0   0.000000
318.000000   1.096758E+0   1.279106E+0   0.000000
319.000000   1.094390E+0   1.281665E+0   0.000000
320.000000   1.091903E+0   1.284302E+0   0.000000
321.000000   1.089308E+0   1.287035E+0   0.000000
322.000000   1.086618E+0   1.289879E+0   0.000000
323.000000   1.083842E+0   1.292850E+0   0.000000
324.000000   1.080992E+0   1.295965E+0   0.000000
325.000000   1.078079E+0   1.299240E+0   0.000000
326.000000   1.075115E+0   1.302690E+0   0.000000
327.000000   1.072110E+0   1.306333E+0   0.000000
328.000000   1.069077E+0   1.310184E+0   0.000000
329.000000   1.066025E+0   1.314258E+0   0.000000
330.000000   1.062967E+0   1.318574E+0   0.000000
331.000000   1.059911E+0   1.323138E+0   0.000000
332.000000   1.056862E+0   1.327932E+0   0.000000
333.000000   1.053822E+0   1.332929E+0   0.000000
334.000000   1.050794E+0   1.338100E+0   0.000000
335.000000   1.047778E+0   1.343419E+0   0.000000
336.000000   1.044779E+0   1.348859E+0   0.000000
337.000000   1.041797E+0   1.354392E+0   0.000000
338.000000   1.038835E+0   1.359991E+0   0.000000
339.000000   1.035895E+0   1.365630E+0   0.000000
340.000000   1.032980E+0   1.371280E+0   0.000000
341.000000   1.030091E+0   1.376915E+0   0.000000
342.000000   1.027231E+0   1.382508E+0   0.000000
343.000000   1.024403E+0   1.388031E+0   0.000000
344.000000   1.021608E+0   1.393457E+0   0.000000
345.000000   1.018849E+0   1.398759E+0   0.000000
346.000000   1.016126E+0   1.403915E+0   0.000000
347.000000   1.013439E+0   1.408931E+0   0.000000
348.000000   1.010785E+0   1.413816E+0   0.000000
349.000000   1.008161E+0   1.418579E+0   0.000000
350.000000   1.005565E+0   1.423232E+0   0.000000
351.000000   1.002994E+0   1.427784E+0   0.000000
352.000000   1.000446E+0   1.432245E+0   0.000000
353.000000   9.979177E-1   1.436625E+0   0.000000
354.000000   9.954073E-1   1.440935E+0   0.000000
355.000000   9.929120E-1   1.445184E+0   0.000000
356.000000   9.904294E-1   1.449383E+0   0.000000
357.000000   9.879568E-1   1.453541E+0   0.000000
358.000000   9.854919E-1   1.457670E+0   0.000000
359.000000   9.830319E-1   1.461778E+0   0.000000
360.000000   9.805745E-1   1.465876E+0   0.000000
Remove Slope = No

Remove Signal Offset = No
Remove Field Offset = No
Cubic Spline Interpolation = No   # Points = 0
Noise Filter = No   Filter Order = 0   Filter Type = Median
Subtract Files = No
[Demagnetizing Field Correction]
Demagnetizing Field Correction = No; Nd = 0.000   (x 4 Pi); Sample Mounted Perpendicular to Field = No
Date and time of last calibration = Friday, June 01, 2018  11:10:26
@@END Instrument Parameters
@@END Parameters
@@Columns
@Column Separator:    
@Column Contents: 
@Number of sections: 7
@Section 0
Column 0: Time since start, Time [s]
Column 1: Raw Temperature, Sample Temperature [degC]
Column 2: Temperature, Sample Temperature [degC]
Column 3: Temperature 2, Sample Temperature [degC]
Column 4: Raw Applied Field, Applied Field [Oe]
Column 5: Applied Field, Applied Field [Oe]
Column 6: Field Angle, Field Angle [deg]
Column 7: Raw Applied Field For Plot , Applied Field [Oe]
Column 8: Applied Field For Plot , Applied Field [Oe]
Column 9: Raw Signal Mx, Moment as measured [memu]
Column 10: Signal X direction, Moment [emu]
@@END Columns
@@End of Header.
Time_since_start   Raw_Temperature   Temperature   Temperature_2   Raw_Applied_Field   Applied_Field   Field_Angle   Raw_Applied_Field_For_Plot_   Applied_Field_For_Plot_   Raw_Signal_Mx   Signal_X_direction      
@Time at start of measurement: 15:52:50
@@Data
New Section: Section 0: 
5.032000E+0   2.231960E+1   2.231960E+1   2.766729E+1   -1.699900E+4   -1.699900E+4   0.000000E+0   -1.699900E+4   -1.699900E+4   1.029519E+0   -1.164803E-5   
1.913300E+1   2.230401E+1   2.230401E+1   2.741641E+1   -1.599900E+4   -1.599900E+4   0.000000E+0   -1.600000E+4   -1.600000E+4   9.656612E-1   -1.548578E-5   
3.271800E+1   2.228231E+1   2.228231E+1   2.728890E+1   -1.499900E+4   -1.499900E+4   0.000000E+0   -1.500000E+4   -1.500000E+4   9.039749E-1   -1.567083E-5   
4.529200E+1   2.228439E+1   2.228439E+1   2.737390E+1   -1.399900E+4   -1.399900E+4   0.000000E+0   -1.400000E+4   -1.400000E+4   8.327377E-1   -2.499161E-5   
5.841800E+1   2.226711E+1   2.226711E+1   2.736129E+1   -1.300000E+4   -1.300000E+4   0.000000E+0   -1.300100E+4   -1.300100E+4   7.667100E-1   -2.916727E-5   
6.996200E+1   2.225991E+1   2.225991E+1   2.733730E+1   -1.199900E+4   -1.199900E+4   0.000000E+0   -1.200100E+4   -1.200100E+4   6.993777E-1   -3.458498E-5   
8.159200E+1   2.225540E+1   2.225540E+1   2.720330E+1   -1.100000E+4   -1.100000E+4   0.000000E+0   -1.100100E+4   -1.100100E+4   6.307433E-1   -4.130423E-5   
9.257500E+1   2.224511E+1   2.224511E+1   2.717101E+1   -9.998000E+3   -9.998000E+3   0.000000E+0   -1.000000E+4   -1.000000E+4   5.651499E-1   -4.492196E-5   
1.028840E+2   2.225039E+1   2.225039E+1   2.733709E+1   -8.999000E+3   -8.999000E+3   0.000000E+0   -9.001000E+3   -9.001000E+3   4.991199E-1   -4.909995E-5   
1.134760E+2   2.224828E+1   2.224828E+1   2.742089E+1   -7.999000E+3   -7.999000E+3   0.000000E+0   -8.000000E+3   -8.000000E+3   4.244043E-1   -6.183570E-5   
1.242630E+2   2.224200E+1   2.224200E+1   2.749828E+1   -7.000000E+3   -7.000000E+3   0.000000E+0   -7.001000E+3   -7.001000E+3   3.614171E-1   -6.297224E-5   
1.346130E+2   2.224789E+1   2.224789E+1   2.771411E+1   -5.999000E+3   -5.999000E+3   0.000000E+0   -6.001000E+3   -6.001000E+3   3.019054E-1   -6.057296E-5   
1.454510E+2   2.225381E+1   2.225381E+1   2.780410E+1   -4.999000E+3   -4.999000E+3   0.000000E+0   -5.001000E+3   -5.001000E+3   2.263201E-1   -7.423986E-5   
1.557600E+2   2.226019E+1   2.226019E+1   2.792059E+1   -3.999000E+3   -3.999000E+3   0.000000E+0   -4.000000E+3   -4.000000E+3   1.598578E-1   -7.872613E-5   
1.660590E+2   2.227529E+1   2.227529E+1   2.775771E+1   -2.999000E+3   -2.999000E+3   0.000000E+0   -3.001000E+3   -3.001000E+3   9.122277E-2   -8.550791E-5   
1.764150E+2   2.228149E+1   2.228149E+1   2.764071E+1   -1.999000E+3   -1.999000E+3   0.000000E+0   -2.001000E+3   -2.001000E+3   3.127652E-2   -8.354300E-5   
1.874740E+2   2.231191E+1   2.231191E+1   2.781249E+1   -1.000000E+3   -1.000000E+3   0.000000E+0   -1.001000E+3   -1.001000E+3   -3.996442E-2   -9.286758E-5   
2.090910E+2   2.232830E+1   2.232830E+1   2.762100E+1   -9.000000E+2   -9.000000E+2   0.000000E+0   -9.020000E+2   -9.020000E+2   -4.821791E-2   -9.499080E-5   
2.168120E+2   2.233700E+1   2.233700E+1   2.775329E+1   -7.990000E+2   -7.990000E+2   0.000000E+0   -8.000000E+2   -8.000000E+2   -5.038989E-2   -9.084965E-5   
2.245740E+2   2.233801E+1   2.233801E+1   2.771420E+1   -7.000000E+2   -7.000000E+2   0.000000E+0   -7.000000E+2   -7.000000E+2   -5.429945E-2   -8.856905E-5   
2.322670E+2   2.234469E+1   2.234469E+1   2.772000E+1   -6.000000E+2   -6.000000E+2   0.000000E+0   -6.000000E+2   -6.000000E+2   -6.472500E-2   -9.280145E-5   
2.400060E+2   2.236151E+1   2.236151E+1   2.774340E+1   -4.990000E+2   -4.990000E+2   0.000000E+0   -5.000000E+2   -5.000000E+2   -6.385616E-2   -8.574465E-5   
2.605460E+2   2.235421E+1   2.235421E+1   2.763830E+1   -4.490000E+2   -4.490000E+2   0.000000E+0   -4.510000E+2   -4.510000E+2   -7.167552E-2   -9.052811E-5   
2.675700E+2   2.236611E+1   2.236611E+1   2.790389E+1   -3.990000E+2   -3.990000E+2   0.000000E+0   -4.000000E+2   -4.000000E+2   -7.124109E-2   -8.693782E-5   
2.746400E+2   2.237161E+1   2.237161E+1   2.782681E+1   -3.490000E+2   -3.490000E+2   0.000000E+0   -3.500000E+2   -3.500000E+2   -8.253529E-2   -9.513265E-5   
2.817000E+2   2.237890E+1   2.237890E+1   2.781521E+1   -2.990000E+2   -2.990000E+2   0.000000E+0   -3.000000E+2   -3.000000E+2   -7.992891E-2   -8.943329E-5   
2.887640E+2   2.238830E+1   2.238830E+1   2.779720E+1   -2.490000E+2   -2.490000E+2   0.000000E+0   -2.500000E+2   -2.500000E+2   -9.078863E-2   -9.719384E-5   
2.958540E+2   2.238729E+1   2.238729E+1   2.767809E+1   -1.990000E+2   -1.990000E+2   0.000000E+0   -2.000000E+2   -2.000000E+2   -8.166638E-2   -8.498159E-5   
3.028540E+2   2.239370E+1   2.239370E+1   2.771761E+1   -1.490000E+2   -1.490000E+2   0.000000E+0   -1.500000E+2   -1.500000E+2   -9.209171E-2   -9.230795E-5   
3.099080E+2   2.239391E+1   2.239391E+1   2.782180E+1   -9.900000E+1   -9.900000E+1   0.000000E+0   -1.000000E+2   -1.000000E+2   -9.382936E-2   -9.095063E-5   
3.318260E+2   2.242581E+1   2.242581E+1   2.795779E+1   -8.900000E+1   -8.900000E+1   0.000000E+0   -9.100000E+1   -9.100000E+1   -9.730453E-2   -9.386725E-5   
3.377500E+2   2.242880E+1   2.242880E+1   2.781271E+1   -7.900000E+1   -7.900000E+1   0.000000E+0   -7.900000E+1   -7.900000E+1   -9.252621E-2   -8.834852E-5   
3.438490E+2   2.243539E+1   2.243539E+1   2.769769E+1   -6.900000E+1   -6.900000E+1   0.000000E+0   -6.900000E+1   -6.900000E+1   -9.904197E-2   -9.424245E-5   
3.497480E+2   2.243911E+1   2.243911E+1   2.761721E+1   -5.900000E+1   -5.900000E+1   0.000000E+0   -5.900000E+1   -5.900000E+1   -9.730453E-2   -9.188697E-5   
3.556050E+2   2.244839E+1   2.244839E+1   2.777169E+1   -4.900000E+1   -4.900000E+1   0.000000E+0   -4.900000E+1   -4.900000E+1   -9.600131E-2   -8.996551E-5   
3.614930E+2   2.244399E+1   2.244399E+1   2.780749E+1   -3.900000E+1   -3.900000E+1   0.000000E+0   -3.900000E+1   -3.900000E+1   -9.687017E-2   -9.021514E-5   
3.673640E+2   2.245410E+1   2.245410E+1   2.772711E+1   -2.900000E+1   -2.900000E+1   0.000000E+0   -2.900000E+1   -2.900000E+1   -9.687010E-2   -8.959623E-5   
3.732080E+2   2.245681E+1   2.245681E+1   2.778329E+1   -1.900000E+1   -1.900000E+1   0.000000E+0   -1.900000E+1   -1.900000E+1   -9.687017E-2   -8.897746E-5   
3.789930E+2   2.246490E+1   2.246490E+1   2.784939E+1   -9.000000E+0   -9.000000E+0   0.000000E+0   -9.000000E+0   -9.000000E+0   -9.773889E-2   -8.922695E-5   
3.847480E+2   2.246230E+1   2.246230E+1   2.783071E+1   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   -9.426380E-2   -8.519650E-5   
3.909170E+2   2.248000E+1   2.248000E+1   2.801461E+1   9.000000E+0   9.000000E+0   0.000000E+0   9.000000E+0   9.000000E+0   -9.817339E-2   -8.854735E-5   
3.972240E+2   2.247851E+1   2.247851E+1   2.806552E+1   1.900000E+1   1.900000E+1   0.000000E+0   1.900000E+1   1.900000E+1   -9.339500E-2   -8.315231E-5   
4.033160E+2   2.248989E+1   2.248989E+1   2.809951E+1   2.900000E+1   2.900000E+1   0.000000E+0   2.900000E+1   2.900000E+1   -9.556695E-2   -8.470442E-5   
4.096320E+2   2.248290E+1   2.248290E+1   2.817901E+1   3.900000E+1   3.900000E+1   0.000000E+0   3.800000E+1   3.800000E+1   -9.556702E-2   -8.414754E-5   
4.163010E+2   2.247949E+1   2.247949E+1   2.792071E+1   4.900000E+1   4.900000E+1   0.000000E+0   4.900000E+1   4.900000E+1   -8.036335E-2   -6.827013E-5   
4.223900E+2   2.248849E+1   2.248849E+1   2.783431E+1   5.900000E+1   5.900000E+1   0.000000E+0   5.900000E+1   5.900000E+1   2.085100E-2   3.351661E-5   
4.287000E+2   2.248531E+1   2.248531E+1   2.779681E+1   6.900000E+1   6.900000E+1   0.000000E+0   6.900000E+1   6.900000E+1   5.082427E-2   6.409497E-5   
4.349680E+2   2.247790E+1   2.247790E+1   2.760009E+1   7.900000E+1   7.900000E+1   0.000000E+0   7.900000E+1   7.900000E+1   5.994654E-2   7.383188E-5   
4.412390E+2   2.248171E+1   2.248171E+1   2.757919E+1   8.900000E+1   8.900000E+1   0.000000E+0   8.900000E+1   8.900000E+1   5.864355E-2   7.314833E-5   
4.475100E+2   2.248409E+1   2.248409E+1   2.768881E+1   9.900000E+1   9.900000E+1   0.000000E+0   9.900000E+1   9.900000E+1   6.429060E-2   7.941163E-5   
4.657970E+2   2.249111E+1   2.249111E+1   2.751739E+1   1.490000E+2   1.490000E+2   0.000000E+0   1.500000E+2   1.500000E+2   5.473381E-2   7.301529E-5   
4.731840E+2   2.248449E+1   2.248449E+1   2.752542E+1   1.990000E+2   1.990000E+2   0.000000E+0   1.980000E+2   1.980000E+2   5.343063E-2   7.468312E-5   
4.805910E+2   2.247411E+1   2.247411E+1   2.750570E+1   2.490000E+2   2.490000E+2   0.000000E+0   2.480000E+2   2.480000E+2   5.125866E-2   7.560633E-5   
4.882220E+2   2.248010E+1   2.248010E+1   2.763220E+1   2.980000E+2   2.980000E+2   0.000000E+0   2.980000E+2   2.980000E+2   4.604595E-2   7.349019E-5   
4.956600E+2   2.246951E+1   2.246951E+1   2.762841E+1   3.480000E+2   3.480000E+2   0.000000E+0   3.480000E+2   3.480000E+2   5.082427E-2   8.136050E-5   
5.030880E+2   2.247189E+1   2.247189E+1   2.773211E+1   3.980000E+2   3.980000E+2   0.000000E+0   3.980000E+2   3.980000E+2   4.474276E-2   7.837597E-5   
5.110170E+2   2.246749E+1   2.246749E+1   2.759249E+1   4.480000E+2   4.480000E+2   0.000000E+0   4.480000E+2   4.480000E+2   4.648034E-2   8.320694E-5   
5.184800E+2   2.245110E+1   2.245110E+1   2.749261E+1   4.980000E+2   4.980000E+2   0.000000E+0   4.980000E+2   4.980000E+2   6.602817E-2   1.058400E-4   
5.394100E+2   2.244891E+1   2.244891E+1   2.757501E+1   5.980000E+2   5.980000E+2   0.000000E+0   6.000000E+2   6.000000E+2   3.214528E-2   7.828477E-5   
5.482000E+2   2.244149E+1   2.244149E+1   2.750060E+1   6.980000E+2   6.980000E+2   0.000000E+0   6.970000E+2   6.970000E+2   2.823572E-2   8.037971E-5   
5.569470E+2   2.243990E+1   2.243990E+1   2.744052E+1   7.980000E+2   7.980000E+2   0.000000E+0   7.970000E+2   7.970000E+2   1.867903E-2   7.701578E-5   
5.662180E+2   2.245519E+1   2.245519E+1   2.770049E+1   8.980000E+2   8.980000E+2   0.000000E+0   8.980000E+2   8.980000E+2   1.781023E-2   8.239763E-5   
5.749630E+2   2.244589E+1   2.244589E+1   2.778591E+1   9.980000E+2   9.980000E+2   0.000000E+0   9.970000E+2   9.970000E+2   1.476946E-2   8.548473E-5   
5.887390E+2   2.243371E+1   2.243371E+1   2.780319E+1   1.999000E+3   1.999000E+3   0.000000E+0   1.998000E+3   1.998000E+3   -5.125868E-2   8.143244E-5   
6.020800E+2   2.242529E+1   2.242529E+1   2.760040E+1   2.999000E+3   2.999000E+3   0.000000E+0   2.998000E+3   2.998000E+3   -1.242370E-1   7.037127E-5   
6.141230E+2   2.242669E+1   2.242669E+1   2.767321E+1   3.999000E+3   3.999000E+3   0.000000E+0   3.998000E+3   3.998000E+3   -1.911340E-1   6.538859E-5   
6.264110E+2   2.240951E+1   2.240951E+1   2.790630E+1   4.998000E+3   4.998000E+3   0.000000E+0   4.998000E+3   4.998000E+3   -2.549898E-1   6.344583E-5   
6.389390E+2   2.240371E+1   2.240371E+1   2.771899E+1   5.999000E+3   5.999000E+3   0.000000E+0   5.998000E+3   5.998000E+3   -3.227563E-1   5.759403E-5   
6.512390E+2   2.239291E+1   2.239291E+1   2.773559E+1   6.998000E+3   6.998000E+3   0.000000E+0   6.997000E+3   6.997000E+3   -3.861778E-1   5.602348E-5   
6.632240E+2   2.240441E+1   2.240441E+1   2.772091E+1   7.999000E+3   7.999000E+3   0.000000E+0   7.998000E+3   7.998000E+3   -4.522055E-1   5.197159E-5   
6.757170E+2   2.238729E+1   2.238729E+1   2.765219E+1   8.998000E+3   8.998000E+3   0.000000E+0   8.998000E+3   8.998000E+3   -5.243149E-1   4.177891E-5   
6.877180E+2   2.239651E+1   2.239651E+1   2.756750E+1   9.999000E+3   9.999000E+3   0.000000E+0   9.998000E+3   9.998000E+3   -5.977293E-1   3.028187E-5   
7.000250E+2   2.239349E+1   2.239349E+1   2.777221E+1   1.099900E+4   1.099900E+4   0.000000E+0   1.099800E+4   1.099800E+4   -6.624539E-1   2.747064E-5   
7.131210E+2   2.238439E+1   2.238439E+1   2.768881E+1   1.199900E+4   1.199900E+4   0.000000E+0   1.199800E+4   1.199800E+4   -7.302193E-1   2.162001E-5   
7.262710E+2   2.238751E+1   2.238751E+1   2.773351E+1   1.299800E+4   1.299800E+4   0.000000E+0   1.299800E+4   1.299800E+4   -7.827813E-1   3.096578E-5   
7.396380E+2   2.238769E+1   2.238769E+1   2.788110E+1   1.399900E+4   1.399900E+4   0.000000E+0   1.399800E+4   1.399800E+4   -8.657512E-1   9.917574E-6   
7.534380E+2   2.238711E+1   2.238711E+1   2.770220E+1   1.499800E+4   1.499800E+4   0.000000E+0   1.499800E+4   1.499800E+4   -9.287377E-1   8.843647E-6   
7.675470E+2   2.238949E+1   2.238949E+1   2.764959E+1   1.599900E+4   1.599900E+4   0.000000E+0   1.599800E+4   1.599800E+4   -9.834699E-1   1.560467E-5   
7.840130E+2   2.236859E+1   2.236859E+1   2.765350E+1   1.699800E+4   1.699800E+4   0.000000E+0   1.699800E+4   1.699800E+4   -1.043853E+0   1.527796E-5   
8.011030E+2   2.236950E+1   2.236950E+1   2.774499E+1   1.600000E+4   1.600000E+4   0.000000E+0   1.600100E+4   1.600100E+4   -9.865104E-1   1.274572E-5   
8.153120E+2   2.236401E+1   2.236401E+1   2.770089E+1   1.499900E+4   1.499900E+4   0.000000E+0   1.500000E+4   1.500000E+4   -9.196118E-1   1.808915E-5   
8.288810E+2   2.236981E+1   2.236981E+1   2.742220E+1   1.400000E+4   1.400000E+4   0.000000E+0   1.400100E+4   1.400100E+4   -8.527205E-1   2.312803E-5   
8.416890E+2   2.237530E+1   2.237530E+1   2.752090E+1   1.299900E+4   1.299900E+4   0.000000E+0   1.300000E+4   1.300000E+4   -7.884280E-1   2.544547E-5   
8.539910E+2   2.236910E+1   2.236910E+1   2.762991E+1   1.199900E+4   1.199900E+4   0.000000E+0   1.200000E+4   1.200000E+4   -7.237027E-1   2.825734E-5   
8.662340E+2   2.236349E+1   2.236349E+1   2.775149E+1   1.099900E+4   1.099900E+4   0.000000E+0   1.100000E+4   1.100000E+4   -6.481190E-1   4.192271E-5   
8.784640E+2   2.235449E+1   2.235449E+1   2.770971E+1   9.999000E+3   9.999000E+3   0.000000E+0   1.000000E+4   1.000000E+4   -5.985980E-1   2.953731E-5   
8.894820E+2   2.234030E+1   2.234030E+1   2.767529E+1   8.999000E+3   8.999000E+3   0.000000E+0   9.000000E+3   9.000000E+3   -5.264869E-1   3.973173E-5   
9.013480E+2   2.233480E+1   2.233480E+1   2.783239E+1   7.999000E+3   7.999000E+3   0.000000E+0   8.000000E+3   8.000000E+3   -4.548120E-1   4.949003E-5   
9.122810E+2   2.234509E+1   2.234509E+1   2.792910E+1   6.998000E+3   6.998000E+3   0.000000E+0   7.000000E+3   7.000000E+3   -3.844401E-1   5.794599E-5   
9.234590E+2   2.234310E+1   2.234310E+1   2.764791E+1   5.999000E+3   5.999000E+3   0.000000E+0   6.000000E+3   6.000000E+3   -3.284036E-1   5.207313E-5   
9.351650E+2   2.233901E+1   2.233901E+1   2.766369E+1   4.998000E+3   4.998000E+3   0.000000E+0   4.999000E+3   4.999000E+3   -2.688909E-1   4.961299E-5   
9.466510E+2   2.232989E+1   2.232989E+1   2.756490E+1   3.999000E+3   3.999000E+3   0.000000E+0   4.000000E+3   4.000000E+3   -1.893965E-1   6.724907E-5   
9.573930E+2   2.232672E+1   2.232672E+1   2.772201E+1   2.999000E+3   2.999000E+3   0.000000E+0   3.001000E+3   3.001000E+3   -1.224995E-1   7.229363E-5   
9.688570E+2   2.233349E+1   2.233349E+1   2.767849E+1   1.999000E+3   1.999000E+3   0.000000E+0   2.000000E+3   2.000000E+3   -5.386503E-2   7.895105E-5   
9.798840E+2   2.233611E+1   2.233611E+1   2.785049E+1   9.990000E+2   9.990000E+2   0.000000E+0   1.000000E+3   1.000000E+3   9.991106E-3   8.089422E-5   
1.002042E+3   2.233441E+1   2.233441E+1   2.767059E+1   8.980000E+2   8.980000E+2   0.000000E+0   9.000000E+2   9.000000E+2   1.303188E-2   7.774523E-5   
1.009966E+3   2.234051E+1   2.234051E+1   2.766189E+1   7.980000E+2   7.980000E+2   0.000000E+0   7.990000E+2   7.990000E+2   1.694144E-2   7.540275E-5   
1.017948E+3   2.234121E+1   2.234121E+1   2.776489E+1   6.980000E+2   6.980000E+2   0.000000E+0   6.990000E+2   6.990000E+2   2.519495E-2   7.746411E-5   
1.025939E+3   2.233499E+1   2.233499E+1   2.768929E+1   5.980000E+2   5.980000E+2   0.000000E+0   5.990000E+2   5.990000E+2   3.692362E-2   8.299903E-5   
1.033848E+3   2.234551E+1   2.234551E+1   2.768170E+1   4.980000E+2   4.980000E+2   0.000000E+0   4.990000E+2   4.990000E+2   3.909563E-2   7.898168E-5   
1.054922E+3   2.235491E+1   2.235491E+1   2.799630E+1   4.490000E+2   4.490000E+2   0.000000E+0   4.500000E+2   4.500000E+2   3.735807E-2   7.421262E-5   
1.062195E+3   2.235311E+1   2.235311E+1   2.790688E+1   3.990000E+2   3.990000E+2   0.000000E+0   3.990000E+2   3.990000E+2   4.908671E-2   8.277981E-5   
1.069838E+3   2.235851E+1   2.235851E+1   2.795599E+1   3.490000E+2   3.490000E+2   0.000000E+0   3.490000E+2   3.490000E+2   4.865231E-2   7.925142E-5   
1.077130E+3   2.236859E+1   2.236859E+1   2.790881E+1   2.980000E+2   2.980000E+2   0.000000E+0   2.990000E+2   2.990000E+2   5.169304E-2   7.919658E-5   
1.084471E+3   2.236630E+1   2.236630E+1   2.770999E+1   2.490000E+2   2.490000E+2   0.000000E+0   2.490000E+2   2.490000E+2   4.995550E-2   7.436565E-5   
1.091763E+3   2.236160E+1   2.236160E+1   2.766140E+1   1.990000E+2   1.990000E+2   0.000000E+0   1.990000E+2   1.990000E+2   5.994654E-2   8.125792E-5   
1.098981E+3   2.237271E+1   2.237271E+1   2.759939E+1   1.490000E+2   1.490000E+2   0.000000E+0   1.490000E+2   1.490000E+2   5.777458E-2   7.599277E-5   
1.106118E+3   2.237219E+1   2.237219E+1   2.767379E+1   9.900000E+1   9.900000E+1   0.000000E+0   9.900000E+1   9.900000E+1   6.559377E-2   8.071419E-5   
1.128600E+3   2.236959E+1   2.236959E+1   2.763879E+1   8.900000E+1   8.900000E+1   0.000000E+0   9.000000E+1   9.000000E+1   6.689693E-2   8.145980E-5   
1.134905E+3   2.237460E+1   2.237460E+1   2.752291E+1   7.900000E+1   7.900000E+1   0.000000E+0   7.900000E+1   7.900000E+1   6.515942E-2   7.904237E-5   
1.141480E+3   2.237209E+1   2.237209E+1   2.758801E+1   6.900000E+1   6.900000E+1   0.000000E+0   6.900000E+1   6.900000E+1   5.647141E-2   6.973951E-5   
1.147703E+3   2.238610E+1   2.238610E+1   2.753039E+1   5.900000E+1   5.900000E+1   0.000000E+0   5.900000E+1   5.900000E+1   6.689705E-2   7.954152E-5   
1.153950E+3   2.238781E+1   2.238781E+1   2.748959E+1   4.900000E+1   4.900000E+1   0.000000E+0   4.900000E+1   4.900000E+1   6.255298E-2   7.458061E-5   
1.160230E+3   2.238671E+1   2.238671E+1   2.763360E+1   3.900000E+1   3.900000E+1   0.000000E+0   3.900000E+1   3.900000E+1   6.429058E-2   7.569858E-5   
1.166498E+3   2.239529E+1   2.239529E+1   2.771029E+1   2.900000E+1   2.900000E+1   0.000000E+0   2.900000E+1   2.900000E+1   6.515942E-2   7.594819E-5   
1.172758E+3   2.238650E+1   2.238650E+1   2.792660E+1   1.900000E+1   1.900000E+1   0.000000E+0   1.900000E+1   1.900000E+1   5.907784E-2   6.925056E-5   
1.178564E+3   2.239099E+1   2.239099E+1   2.809121E+1   9.000000E+0   9.000000E+0   0.000000E+0   9.000000E+0   9.000000E+0   6.515942E-2   7.471051E-5   
1.184248E+3   2.239391E+1   2.239391E+1   2.792169E+1   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   6.602823E-2   7.502197E-5   
1.190074E+3   2.239001E+1   2.239001E+1   2.778790E+1   -9.000000E+0   -9.000000E+0   0.000000E+0   -9.000000E+0   -9.000000E+0   6.255298E-2   7.099136E-5   
1.195980E+3   2.238070E+1   2.238070E+1   2.794430E+1   -1.900000E+1   -1.900000E+1   0.000000E+0   -1.900000E+1   -1.900000E+1   5.994656E-2   6.776730E-5   
1.201915E+3   2.239059E+1   2.239059E+1   2.803411E+1   -2.900000E+1   -2.900000E+1   0.000000E+0   -2.800000E+1   -2.800000E+1   6.689705E-2   7.415765E-5   
1.207799E+3   2.239370E+1   2.239370E+1   2.805041E+1   -3.900000E+1   -3.900000E+1   0.000000E+0   -3.900000E+1   -3.900000E+1   6.602825E-2   7.260853E-5   
1.213706E+3   2.240301E+1   2.240301E+1   2.791021E+1   -4.900000E+1   -4.900000E+1   0.000000E+0   -4.900000E+1   -4.900000E+1   6.602819E-2   7.198964E-5   
1.219637E+3   2.239459E+1   2.239459E+1   2.777169E+1   -5.900000E+1   -5.900000E+1   0.000000E+0   -5.900000E+1   -5.900000E+1   -2.171980E-2   -1.633693E-5   
1.225499E+3   2.240740E+1   2.240740E+1   2.766180E+1   -6.900000E+1   -6.900000E+1   0.000000E+0   -6.900000E+1   -6.900000E+1   -7.645370E-2   -7.166455E-5   
1.231380E+3   2.239871E+1   2.239871E+1   2.765710E+1   -7.900000E+1   -7.900000E+1   0.000000E+0   -7.800000E+1   -7.800000E+1   -9.035434E-2   -8.611576E-5   
1.237258E+3   2.240521E+1   2.240521E+1   2.764211E+1   -8.900000E+1   -8.900000E+1   0.000000E+0   -8.900000E+1   -8.900000E+1   -9.296072E-2   -8.940166E-5   
1.243258E+3   2.240841E+1   2.240841E+1   2.769540E+1   -9.900000E+1   -9.900000E+1   0.000000E+0   -9.900000E+1   -9.900000E+1   -7.906004E-2   -7.612620E-5   
1.260626E+3   2.240820E+1   2.240820E+1   2.766009E+1   -1.500000E+2   -1.500000E+2   0.000000E+0   -1.520000E+2   -1.520000E+2   -8.687918E-2   -8.722158E-5   
1.267805E+3   2.241830E+1   2.241830E+1   2.763021E+1   -1.990000E+2   -1.990000E+2   0.000000E+0   -1.980000E+2   -1.980000E+2   -9.122313E-2   -9.441019E-5   
1.274984E+3   2.242031E+1   2.242031E+1   2.740811E+1   -2.490000E+2   -2.490000E+2   0.000000E+0   -2.480000E+2   -2.480000E+2   -7.645370E-2   -8.274172E-5   
1.282363E+3   2.241299E+1   2.241299E+1   2.735729E+1   -2.990000E+2   -2.990000E+2   0.000000E+0   -2.980000E+2   -2.980000E+2   -8.253523E-2   -9.191464E-5   
1.289553E+3   2.241519E+1   2.241519E+1   2.734680E+1   -3.490000E+2   -3.490000E+2   0.000000E+0   -3.480000E+2   -3.480000E+2   -7.558490E-2   -8.806169E-5   
1.296725E+3   2.241549E+1   2.241549E+1   2.756149E+1   -3.990000E+2   -3.990000E+2   0.000000E+0   -3.980000E+2   -3.980000E+2   -7.819133E-2   -9.376110E-5   
1.303930E+3   2.242239E+1   2.242239E+1   2.749911E+1   -4.490000E+2   -4.490000E+2   0.000000E+0   -4.480000E+2   -4.480000E+2   -7.124093E-2   -8.990808E-5   
1.311077E+3   2.242300E+1   2.242300E+1   2.750939E+1   -4.990000E+2   -4.990000E+2   0.000000E+0   -4.980000E+2   -4.980000E+2   -7.297859E-2   -9.473912E-5   
1.331375E+3   2.241619E+1   2.241619E+1   2.773651E+1   -6.000000E+2   -6.000000E+2   0.000000E+0   -6.020000E+2   -6.020000E+2   -6.689701E-2   -9.509623E-5   
1.339125E+3   2.241940E+1   2.241940E+1   2.769161E+1   -6.990000E+2   -6.990000E+2   0.000000E+0   -6.980000E+2   -6.980000E+2   -5.038991E-2   -8.453753E-5   
1.346981E+3   2.241119E+1   2.241119E+1   2.773150E+1   -7.990000E+2   -7.990000E+2   0.000000E+0   -7.980000E+2   -7.980000E+2   -5.473381E-2   -9.506781E-5   
1.355016E+3   2.240801E+1   2.240801E+1   2.772579E+1   -8.990000E+2   -8.990000E+2   0.000000E+0   -8.980000E+2   -8.980000E+2   -4.604594E-2   -9.257229E-5   
1.362872E+3   2.241079E+1   2.241079E+1   2.776510E+1   -9.990000E+2   -9.990000E+2   0.000000E+0   -9.980000E+2   -9.980000E+2   -3.648931E-2   -8.920842E-5   
1.377182E+3   2.240551E+1   2.240551E+1   2.776101E+1   -1.998000E+3   -1.998000E+3   0.000000E+0   -1.997000E+3   -1.997000E+3   1.911343E-2   -9.545296E-5   
1.389958E+3   2.241921E+1   2.241921E+1   2.791461E+1   -2.998000E+3   -2.998000E+3   0.000000E+0   -2.998000E+3   -2.998000E+3   9.382951E-2   -8.271672E-5   
1.401760E+3   2.240429E+1   2.240429E+1   2.796569E+1   -3.998000E+3   -3.998000E+3   0.000000E+0   -3.997000E+3   -3.997000E+3   1.589889E-1   -7.940902E-5   
1.413043E+3   2.241589E+1   2.241589E+1   2.764889E+1   -4.999000E+3   -4.999000E+3   0.000000E+0   -4.998000E+3   -4.998000E+3   2.145916E-1   -8.577740E-5   
1.425392E+3   2.240829E+1   2.240829E+1   2.762530E+1   -5.999000E+3   -5.999000E+3   0.000000E+0   -5.998000E+3   -5.998000E+3   2.901769E-1   -7.211043E-5   
1.436327E+3   2.240890E+1   2.240890E+1   2.775491E+1   -6.999000E+3   -6.999000E+3   0.000000E+0   -6.997000E+3   -6.997000E+3   3.640237E-1   -6.011923E-5   
1.448125E+3   2.242739E+1   2.242739E+1   2.773931E+1   -7.998000E+3   -7.998000E+3   0.000000E+0   -7.997000E+3   -7.997000E+3   4.248385E-1   -6.121603E-5   
1.460740E+3   2.243041E+1   2.243041E+1   2.782849E+1   -8.999000E+3   -8.999000E+3   0.000000E+0   -8.998000E+3   -8.998000E+3   5.030297E-1   -4.500627E-5   
1.472591E+3   2.241851E+1   2.241851E+1   2.758560E+1   -9.998000E+3   -9.998000E+3   0.000000E+0   -9.997000E+3   -9.997000E+3   5.568958E-1   -5.298666E-5   
1.484207E+3   2.241619E+1   2.241619E+1   2.757781E+1   -1.099900E+4   -1.099900E+4   0.000000E+0   -1.099800E+4   -1.099800E+4   6.281372E-1   -4.372354E-5   
1.497382E+3   2.240341E+1   2.240341E+1   2.770349E+1   -1.199900E+4   -1.199900E+4   0.000000E+0   -1.199800E+4   -1.199800E+4   6.932958E-1   -4.047845E-5   
1.509476E+3   2.239929E+1   2.239929E+1   2.755139E+1   -1.299900E+4   -1.299900E+4   0.000000E+0   -1.299800E+4   -1.299800E+4   7.654069E-1   -3.028410E-5   
1.522585E+3   2.238830E+1   2.238830E+1   2.770779E+1   -1.399800E+4   -1.399800E+4   0.000000E+0   -1.399700E+4   -1.399700E+4   8.340423E-1   -2.350202E-5   
1.535674E+3   2.237469E+1   2.237469E+1   2.784081E+1   -1.499800E+4   -1.499800E+4   0.000000E+0   -1.499700E+4   -1.499700E+4   9.078841E-1   -1.157773E-5   
1.550305E+3   2.236669E+1   2.236669E+1   2.793401E+1   -1.599800E+4   -1.599800E+4   0.000000E+0   -1.599700E+4   -1.599700E+4   9.634894E-1   -1.747572E-5   
1.565940E+3   2.237780E+1   2.237780E+1   2.763329E+1   -1.699900E+4   -1.699900E+4   0.000000E+0   -1.699800E+4   -1.699800E+4   1.028649E+0   -1.246000E-5   
@@END Data.
@Time at end of measurement: 16:19:01
@Instrument  Changes:
@Emu Range: 2 mV
@END Instrument  Changes:
@@Final Manipulated Data
New Section: Section 0: 
5.032000E+0   2.231960E+1   2.231960E+1   2.766729E+1   -1.699900E+4   -1.699900E+4   0.000000E+0   -1.699900E+4   -1.699900E+4   1.029519E+0   -1.164803E-5   
1.913300E+1   2.230401E+1   2.230401E+1   2.741641E+1   -1.599900E+4   -1.599900E+4   0.000000E+0   -1.600000E+4   -1.600000E+4   9.656612E-1   -1.548578E-5   
3.271800E+1   2.228231E+1   2.228231E+1   2.728890E+1   -1.499900E+4   -1.499900E+4   0.000000E+0   -1.500000E+4   -1.500000E+4   9.039749E-1   -1.567083E-5   
4.529200E+1   2.228439E+1   2.228439E+1   2.737390E+1   -1.399900E+4   -1.399900E+4   0.000000E+0   -1.400000E+4   -1.400000E+4   8.327377E-1   -2.499161E-5   
5.841800E+1   2.226711E+1   2.226711E+1   2.736129E+1   -1.300000E+4   -1.300000E+4   0.000000E+0   -1.300100E+4   -1.300100E+4   7.667100E-1   -2.916727E-5   
6.996200E+1   2.225991E+1   2.225991E+1   2.733730E+1   -1.199900E+4   -1.199900E+4   0.000000E+0   -1.200100E+4   -1.200100E+4   6.993777E-1   -3.458498E-5   
8.159200E+1   2.225540E+1   2.225540E+1   2.720330E+1   -1.100000E+4   -1.100000E+4   0.000000E+0   -1.100100E+4   -1.100100E+4   6.307433E-1   -4.130423E-5   
9.257500E+1   2.224511E+1   2.224511E+1   2.717101E+1   -9.998000E+3   -9.998000E+3   0.000000E+0   -1.000000E+4   -1.000000E+4   5.651499E-1   -4.492196E-5   
1.028840E+2   2.225039E+1   2.225039E+1   2.733709E+1   -8.999000E+3   -8.999000E+3   0.000000E+0   -9.001000E+3   -9.001000E+3   4.991199E-1   -4.909995E-5   
1.134760E+2   2.224828E+1   2.224828E+1   2.742089E+1   -7.999000E+3   -7.999000E+3   0.000000E+0   -8.000000E+3   -8.000000E+3   4.244043E-1   -6.183570E-5   
1.242630E+2   2.224200E+1   2.224200E+1   2.749828E+1   -7.000000E+3   -7.000000E+3   0.000000E+0   -7.001000E+3   -7.001000E+3   3.614171E-1   -6.297224E-5   
1.346130E+2   2.224789E+1   2.224789E+1   2.771411E+1   -5.999000E+3   -5.999000E+3   0.000000E+0   -6.001000E+3   -6.001000E+3   3.019054E-1   -6.057296E-5   
1.454510E+2   2.225381E+1   2.225381E+1   2.780410E+1   -4.999000E+3   -4.999000E+3   0.000000E+0   -5.001000E+3   -5.001000E+3   2.263201E-1   -7.423986E-5   
1.557600E+2   2.226019E+1   2.226019E+1   2.792059E+1   -3.999000E+3   -3.999000E+3   0.000000E+0   -4.000000E+3   -4.000000E+3   1.598578E-1   -7.872613E-5   
1.660590E+2   2.227529E+1   2.227529E+1   2.775771E+1   -2.999000E+3   -2.999000E+3   0.000000E+0   -3.001000E+3   -3.001000E+3   9.122277E-2   -8.550791E-5   
1.764150E+2   2.228149E+1   2.228149E+1   2.764071E+1   -1.999000E+3   -1.999000E+3   0.000000E+0   -2.001000E+3   -2.001000E+3   3.127652E-2   -8.354300E-5   
1.874740E+2   2.231191E+1   2.231191E+1   2.781249E+1   -1.000000E+3   -1.000000E+3   0.000000E+0   -1.001000E+3   -1.001000E+3   -3.996442E-2   -9.286758E-5   
2.090910E+2   2.232830E+1   2.232830E+1   2.762100E+1   -9.000000E+2   -9.000000E+2   0.000000E+0   -9.020000E+2   -9.020000E+2   -4.821791E-2   -9.499080E-5   
2.168120E+2   2.233700E+1   2.233700E+1   2.775329E+1   -7.990000E+2   -7.990000E+2   0.000000E+0   -8.000000E+2   -8.000000E+2   -5.038989E-2   -9.084965E-5   
2.245740E+2   2.233801E+1   2.233801E+1   2.771420E+1   -7.000000E+2   -7.000000E+2   0.000000E+0   -7.000000E+2   -7.000000E+2   -5.429945E-2   -8.856905E-5   
2.322670E+2   2.234469E+1   2.234469E+1   2.772000E+1   -6.000000E+2   -6.000000E+2   0.000000E+0   -6.000000E+2   -6.000000E+2   -6.472500E-2   -9.280145E-5   
2.400060E+2   2.236151E+1   2.236151E+1   2.774340E+1   -4.990000E+2   -4.990000E+2   0.000000E+0   -5.000000E+2   -5.000000E+2   -6.385616E-2   -8.574465E-5   
2.605460E+2   2.235421E+1   2.235421E+1   2.763830E+1   -4.490000E+2   -4.490000E+2   0.000000E+0   -4.510000E+2   -4.510000E+2   -7.167552E-2   -9.052811E-5   
2.675700E+2   2.236611E+1   2.236611E+1   2.790389E+1   -3.990000E+2   -3.990000E+2   0.000000E+0   -4.000000E+2   -4.000000E+2   -7.124109E-2   -8.693782E-5   
2.746400E+2   2.237161E+1   2.237161E+1   2.782681E+1   -3.490000E+2   -3.490000E+2   0.000000E+0   -3.500000E+2   -3.500000E+2   -8.253529E-2   -9.513265E-5   
2.817000E+2   2.237890E+1   2.237890E+1   2.781521E+1   -2.990000E+2   -2.990000E+2   0.000000E+0   -3.000000E+2   -3.000000E+2   -7.992891E-2   -8.943329E-5   
2.887640E+2   2.238830E+1   2.238830E+1   2.779720E+1   -2.490000E+2   -2.490000E+2   0.000000E+0   -2.500000E+2   -2.500000E+2   -9.078863E-2   -9.719384E-5   
2.958540E+2   2.238729E+1   2.238729E+1   2.767809E+1   -1.990000E+2   -1.990000E+2   0.000000E+0   -2.000000E+2   -2.000000E+2   -8.166638E-2   -8.498159E-5   
3.028540E+2   2.239370E+1   2.239370E+1   2.771761E+1   -1.490000E+2   -1.490000E+2   0.000000E+0   -1.500000E+2   -1.500000E+2   -9.209171E-2   -9.230795E-5   
3.099080E+2   2.239391E+1   2.239391E+1   2.782180E+1   -9.900000E+1   -9.900000E+1   0.000000E+0   -1.000000E+2   -1.000000E+2   -9.382936E-2   -9.095063E-5   
3.318260E+2   2.242581E+1   2.242581E+1   2.795779E+1   -8.900000E+1   -8.900000E+1   0.000000E+0   -9.100000E+1   -9.100000E+1   -9.730453E-2   -9.386725E-5   
3.377500E+2   2.242880E+1   2.242880E+1   2.781271E+1   -7.900000E+1   -7.900000E+1   0.000000E+0   -7.900000E+1   -7.900000E+1   -9.252621E-2   -8.834852E-5   
3.438490E+2   2.243539E+1   2.243539E+1   2.769769E+1   -6.900000E+1   -6.900000E+1   0.000000E+0   -6.900000E+1   -6.900000E+1   -9.904197E-2   -9.424245E-5   
3.497480E+2   2.243911E+1   2.243911E+1   2.761721E+1   -5.900000E+1   -5.900000E+1   0.000000E+0   -5.900000E+1   -5.900000E+1   -9.730453E-2   -9.188697E-5   
3.556050E+2   2.244839E+1   2.244839E+1   2.777169E+1   -4.900000E+1   -4.900000E+1   0.000000E+0   -4.900000E+1   -4.900000E+1   -9.600131E-2   -8.996551E-5   
3.614930E+2   2.244399E+1   2.244399E+1   2.780749E+1   -3.900000E+1   -3.900000E+1   0.000000E+0   -3.900000E+1   -3.900000E+1   -9.687017E-2   -9.021514E-5   
3.673640E+2   2.245410E+1   2.245410E+1   2.772711E+1   -2.900000E+1   -2.900000E+1   0.000000E+0   -2.900000E+1   -2.900000E+1   -9.687010E-2   -8.959623E-5   
3.732080E+2   2.245681E+1   2.245681E+1   2.778329E+1   -1.900000E+1   -1.900000E+1   0.000000E+0   -1.900000E+1   -1.900000E+1   -9.687017E-2   -8.897746E-5   
3.789930E+2   2.246490E+1   2.246490E+1   2.784939E+1   -9.000000E+0   -9.000000E+0   0.000000E+0   -9.000000E+0   -9.000000E+0   -9.773889E-2   -8.922695E-5   
3.847480E+2   2.246230E+1   2.246230E+1   2.783071E+1   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   -9.426380E-2   -8.519650E-5   
3.909170E+2   2.248000E+1   2.248000E+1   2.801461E+1   9.000000E+0   9.000000E+0   0.000000E+0   9.000000E+0   9.000000E+0   -9.817339E-2   -8.854735E-5   
3.972240E+2   2.247851E+1   2.247851E+1   2.806552E+1   1.900000E+1   1.900000E+1   0.000000E+0   1.900000E+1   1.900000E+1   -9.339500E-2   -8.315231E-5   
4.033160E+2   2.248989E+1   2.248989E+1   2.809951E+1   2.900000E+1   2.900000E+1   0.000000E+0   2.900000E+1   2.900000E+1   -9.556695E-2   -8.470442E-5   
4.096320E+2   2.248290E+1   2.248290E+1   2.817901E+1   3.900000E+1   3.900000E+1   0.000000E+0   3.800000E+1   3.800000E+1   -9.556702E-2   -8.414754E-5   
4.163010E+2   2.247949E+1   2.247949E+1   2.792071E+1   4.900000E+1   4.900000E+1   0.000000E+0   4.900000E+1   4.900000E+1   -8.036335E-2   -6.827013E-5   
4.223900E+2   2.248849E+1   2.248849E+1   2.783431E+1   5.900000E+1   5.900000E+1   0.000000E+0   5.900000E+1   5.900000E+1   2.085100E-2   3.351661E-5   
4.287000E+2   2.248531E+1   2.248531E+1   2.779681E+1   6.900000E+1   6.900000E+1   0.000000E+0   6.900000E+1   6.900000E+1   5.082427E-2   6.409497E-5   
4.349680E+2   2.247790E+1   2.247790E+1   2.760009E+1   7.900000E+1   7.900000E+1   0.000000E+0   7.900000E+1   7.900000E+1   5.994654E-2   7.383188E-5   
4.412390E+2   2.248171E+1   2.248171E+1   2.757919E+1   8.900000E+1   8.900000E+1   0.000000E+0   8.900000E+1   8.900000E+1   5.864355E-2   7.314833E-5   
4.475100E+2   2.248409E+1   2.248409E+1   2.768881E+1   9.900000E+1   9.900000E+1   0.000000E+0   9.900000E+1   9.900000E+1   6.429060E-2   7.941163E-5   
4.657970E+2   2.249111E+1   2.249111E+1   2.751739E+1   1.490000E+2   1.490000E+2   0.000000E+0   1.500000E+2   1.500000E+2   5.473381E-2   7.301529E-5   
4.731840E+2   2.248449E+1   2.248449E+1   2.752542E+1   1.990000E+2   1.990000E+2   0.000000E+0   1.980000E+2   1.980000E+2   5.343063E-2   7.468312E-5   
4.805910E+2   2.247411E+1   2.247411E+1   2.750570E+1   2.490000E+2   2.490000E+2   0.000000E+0   2.480000E+2   2.480000E+2   5.125866E-2   7.560633E-5   
4.882220E+2   2.248010E+1   2.248010E+1   2.763220E+1   2.980000E+2   2.980000E+2   0.000000E+0   2.980000E+2   2.980000E+2   4.604595E-2   7.349019E-5   
4.956600E+2   2.246951E+1   2.246951E+1   2.762841E+1   3.480000E+2   3.480000E+2   0.000000E+0   3.480000E+2   3.480000E+2   5.082427E-2   8.136050E-5   
5.030880E+2   2.247189E+1   2.247189E+1   2.773211E+1   3.980000E+2   3.980000E+2   0.000000E+0   3.980000E+2   3.980000E+2   4.474276E-2   7.837597E-5   
5.110170E+2   2.246749E+1   2.246749E+1   2.759249E+1   4.480000E+2   4.480000E+2   0.000000E+0   4.480000E+2   4.480000E+2   4.648034E-2   8.320694E-5   
5.184800E+2   2.245110E+1   2.245110E+1   2.749261E+1   4.980000E+2   4.980000E+2   0.000000E+0   4.980000E+2   4.980000E+2   6.602817E-2   1.058400E-4   
5.394100E+2   2.244891E+1   2.244891E+1   2.757501E+1   5.980000E+2   5.980000E+2   0.000000E+0   6.000000E+2   6.000000E+2   3.214528E-2   7.828477E-5   
5.482000E+2   2.244149E+1   2.244149E+1   2.750060E+1   6.980000E+2   6.980000E+2   0.000000E+0   6.970000E+2   6.970000E+2   2.823572E-2   8.037971E-5   
5.569470E+2   2.243990E+1   2.243990E+1   2.744052E+1   7.980000E+2   7.980000E+2   0.000000E+0   7.970000E+2   7.970000E+2   1.867903E-2   7.701578E-5   
5.662180E+2   2.245519E+1   2.245519E+1   2.770049E+1   8.980000E+2   8.980000E+2   0.000000E+0   8.980000E+2   8.980000E+2   1.781023E-2   8.239763E-5   
5.749630E+2   2.244589E+1   2.244589E+1   2.778591E+1   9.980000E+2   9.980000E+2   0.000000E+0   9.970000E+2   9.970000E+2   1.476946E-2   8.548473E-5   
5.887390E+2   2.243371E+1   2.243371E+1   2.780319E+1   1.999000E+3   1.999000E+3   0.000000E+0   1.998000E+3   1.998000E+3   -5.125868E-2   8.143244E-5   
6.020800E+2   2.242529E+1   2.242529E+1   2.760040E+1   2.999000E+3   2.999000E+3   0.000000E+0   2.998000E+3   2.998000E+3   -1.242370E-1   7.037127E-5   
6.141230E+2   2.242669E+1   2.242669E+1   2.767321E+1   3.999000E+3   3.999000E+3   0.000000E+0   3.998000E+3   3.998000E+3   -1.911340E-1   6.538859E-5   
6.264110E+2   2.240951E+1   2.240951E+1   2.790630E+1   4.998000E+3   4.998000E+3   0.000000E+0   4.998000E+3   4.998000E+3   -2.549898E-1   6.344583E-5   
6.389390E+2   2.240371E+1   2.240371E+1   2.771899E+1   5.999000E+3   5.999000E+3   0.000000E+0   5.998000E+3   5.998000E+3   -3.227563E-1   5.759403E-5   
6.512390E+2   2.239291E+1   2.239291E+1   2.773559E+1   6.998000E+3   6.998000E+3   0.000000E+0   6.997000E+3   6.997000E+3   -3.861778E-1   5.602348E-5   
6.632240E+2   2.240441E+1   2.240441E+1   2.772091E+1   7.999000E+3   7.999000E+3   0.000000E+0   7.998000E+3   7.998000E+3   -4.522055E-1   5.197159E-5   
6.757170E+2   2.238729E+1   2.238729E+1   2.765219E+1   8.998000E+3   8.998000E+3   0.000000E+0   8.998000E+3   8.998000E+3   -5.243149E-1   4.177891E-5   
6.877180E+2   2.239651E+1   2.239651E+1   2.756750E+1   9.999000E+3   9.999000E+3   0.000000E+0   9.998000E+3   9.998000E+3   -5.977293E-1   3.028187E-5   
7.000250E+2   2.239349E+1   2.239349E+1   2.777221E+1   1.099900E+4   1.099900E+4   0.000000E+0   1.099800E+4   1.099800E+4   -6.624539E-1   2.747064E-5   
7.131210E+2   2.238439E+1   2.238439E+1   2.768881E+1   1.199900E+4   1.199900E+4   0.000000E+0   1.199800E+4   1.199800E+4   -7.302193E-1   2.162001E-5   
7.262710E+2   2.238751E+1   2.238751E+1   2.773351E+1   1.299800E+4   1.299800E+4   0.000000E+0   1.299800E+4   1.299800E+4   -7.827813E-1   3.096578E-5   
7.396380E+2   2.238769E+1   2.238769E+1   2.788110E+1   1.399900E+4   1.399900E+4   0.000000E+0   1.399800E+4   1.399800E+4   -8.657512E-1   9.917574E-6   
7.534380E+2   2.238711E+1   2.238711E+1   2.770220E+1   1.499800E+4   1.499800E+4   0.000000E+0   1.499800E+4   1.499800E+4   -9.287377E-1   8.843647E-6   
7.675470E+2   2.238949E+1   2.238949E+1   2.764959E+1   1.599900E+4   1.599900E+4   0.000000E+0   1.599800E+4   1.599800E+4   -9.834699E-1   1.560467E-5   
7.840130E+2   2.236859E+1   2.236859E+1   2.765350E+1   1.699800E+4   1.699800E+4   0.000000E+0   1.699800E+4   1.699800E+4   -1.043853E+0   1.527796E-5   
8.011030E+2   2.236950E+1   2.236950E+1   2.774499E+1   1.600000E+4   1.600000E+4   0.000000E+0   1.600100E+4   1.600100E+4   -9.865104E-1   1.274572E-5   
8.153120E+2   2.236401E+1   2.236401E+1   2.770089E+1   1.499900E+4   1.499900E+4   0.000000E+0   1.500000E+4   1.500000E+4   -9.196118E-1   1.808915E-5   
8.288810E+2   2.236981E+1   2.236981E+1   2.742220E+1   1.400000E+4   1.400000E+4   0.000000E+0   1.400100E+4   1.400100E+4   -8.527205E-1   2.312803E-5   
8.416890E+2   2.237530E+1   2.237530E+1   2.752090E+1   1.299900E+4   1.299900E+4   0.000000E+0   1.300000E+4   1.300000E+4   -7.884280E-1   2.544547E-5   
8.539910E+2   2.236910E+1   2.236910E+1   2.762991E+1   1.199900E+4   1.199900E+4   0.000000E+0   1.200000E+4   1.200000E+4   -7.237027E-1   2.825734E-5   
8.662340E+2   2.236349E+1   2.236349E+1   2.775149E+1   1.099900E+4   1.099900E+4   0.000000E+0   1.100000E+4   1.100000E+4   -6.481190E-1   4.192271E-5   
8.784640E+2   2.235449E+1   2.235449E+1   2.770971E+1   9.999000E+3   9.999000E+3   0.000000E+0   1.000000E+4   1.000000E+4   -5.985980E-1   2.953731E-5   
8.894820E+2   2.234030E+1   2.234030E+1   2.767529E+1   8.999000E+3   8.999000E+3   0.000000E+0   9.000000E+3   9.000000E+3   -5.264869E-1   3.973173E-5   
9.013480E+2   2.233480E+1   2.233480E+1   2.783239E+1   7.999000E+3   7.999000E+3   0.000000E+0   8.000000E+3   8.000000E+3   -4.548120E-1   4.949003E-5   
9.122810E+2   2.234509E+1   2.234509E+1   2.792910E+1   6.998000E+3   6.998000E+3   0.000000E+0   7.000000E+3   7.000000E+3   -3.844401E-1   5.794599E-5   
9.234590E+2   2.234310E+1   2.234310E+1   2.764791E+1   5.999000E+3   5.999000E+3   0.000000E+0   6.000000E+3   6.000000E+3   -3.284036E-1   5.207313E-5   
9.351650E+2   2.233901E+1   2.233901E+1   2.766369E+1   4.998000E+3   4.998000E+3   0.000000E+0   4.999000E+3   4.999000E+3   -2.688909E-1   4.961299E-5   
9.466510E+2   2.232989E+1   2.232989E+1   2.756490E+1   3.999000E+3   3.999000E+3   0.000000E+0   4.000000E+3   4.000000E+3   -1.893965E-1   6.724907E-5   
9.573930E+2   2.232672E+1   2.232672E+1   2.772201E+1   2.999000E+3   2.999000E+3   0.000000E+0   3.001000E+3   3.001000E+3   -1.224995E-1   7.229363E-5   
9.688570E+2   2.233349E+1   2.233349E+1   2.767849E+1   1.999000E+3   1.999000E+3   0.000000E+0   2.000000E+3   2.000000E+3   -5.386503E-2   7.895105E-5   
9.798840E+2   2.233611E+1   2.233611E+1   2.785049E+1   9.990000E+2   9.990000E+2   0.000000E+0   1.000000E+3   1.000000E+3   9.991106E-3   8.089422E-5   
1.002042E+3   2.233441E+1   2.233441E+1   2.767059E+1   8.980000E+2   8.980000E+2   0.000000E+0   9.000000E+2   9.000000E+2   1.303188E-2   7.774523E-5   
1.009966E+3   2.234051E+1   2.234051E+1   2.766189E+1   7.980000E+2   7.980000E+2   0.000000E+0   7.990000E+2   7.990000E+2   1.694144E-2   7.540275E-5   
1.017948E+3   2.234121E+1   2.234121E+1   2.776489E+1   6.980000E+2   6.980000E+2   0.000000E+0   6.990000E+2   6.990000E+2   2.519495E-2   7.746411E-5   
1.025939E+3   2.233499E+1   2.233499E+1   2.768929E+1   5.980000E+2   5.980000E+2   0.000000E+0   5.990000E+2   5.990000E+2   3.692362E-2   8.299903E-5   
1.033848E+3   2.234551E+1   2.234551E+1   2.768170E+1   4.980000E+2   4.980000E+2   0.000000E+0   4.990000E+2   4.990000E+2   3.909563E-2   7.898168E-5   
1.054922E+3   2.235491E+1   2.235491E+1   2.799630E+1   4.490000E+2   4.490000E+2   0.000000E+0   4.500000E+2   4.500000E+2   3.735807E-2   7.421262E-5   
1.062195E+3   2.235311E+1   2.235311E+1   2.790688E+1   3.990000E+2   3.990000E+2   0.000000E+0   3.990000E+2   3.990000E+2   4.908671E-2   8.277981E-5   
1.069838E+3   2.235851E+1   2.235851E+1   2.795599E+1   3.490000E+2   3.490000E+2   0.000000E+0   3.490000E+2   3.490000E+2   4.865231E-2   7.925142E-5   
1.077130E+3   2.236859E+1   2.236859E+1   2.790881E+1   2.980000E+2   2.980000E+2   0.000000E+0   2.990000E+2   2.990000E+2   5.169304E-2   7.919658E-5   
1.084471E+3   2.236630E+1   2.236630E+1   2.770999E+1   2.490000E+2   2.490000E+2   0.000000E+0   2.490000E+2   2.490000E+2   4.995550E-2   7.436565E-5   
1.091763E+3   2.236160E+1   2.236160E+1   2.766140E+1   1.990000E+2   1.990000E+2   0.000000E+0   1.990000E+2   1.990000E+2   5.994654E-2   8.125792E-5   
1.098981E+3   2.237271E+1   2.237271E+1   2.759939E+1   1.490000E+2   1.490000E+2   0.000000E+0   1.490000E+2   1.490000E+2   5.777458E-2   7.599277E-5   
1.106118E+3   2.237219E+1   2.237219E+1   2.767379E+1   9.900000E+1   9.900000E+1   0.000000E+0   9.900000E+1   9.900000E+1   6.559377E-2   8.071419E-5   
1.128600E+3   2.236959E+1   2.236959E+1   2.763879E+1   8.900000E+1   8.900000E+1   0.000000E+0   9.000000E+1   9.000000E+1   6.689693E-2   8.145980E-5   
1.134905E+3   2.237460E+1   2.237460E+1   2.752291E+1   7.900000E+1   7.900000E+1   0.000000E+0   7.900000E+1   7.900000E+1   6.515942E-2   7.904237E-5   
1.141480E+3   2.237209E+1   2.237209E+1   2.758801E+1   6.900000E+1   6.900000E+1   0.000000E+0   6.900000E+1   6.900000E+1   5.647141E-2   6.973951E-5   
1.147703E+3   2.238610E+1   2.238610E+1   2.753039E+1   5.900000E+1   5.900000E+1   0.000000E+0   5.900000E+1   5.900000E+1   6.689705E-2   7.954152E-5   
1.153950E+3   2.238781E+1   2.238781E+1   2.748959E+1   4.900000E+1   4.900000E+1   0.000000E+0   4.900000E+1   4.900000E+1   6.255298E-2   7.458061E-5   
1.160230E+3   2.238671E+1   2.238671E+1   2.763360E+1   3.900000E+1   3.900000E+1   0.000000E+0   3.900000E+1   3.900000E+1   6.429058E-2   7.569858E-5   
1.166498E+3   2.239529E+1   2.239529E+1   2.771029E+1   2.900000E+1   2.900000E+1   0.000000E+0   2.900000E+1   2.900000E+1   6.515942E-2   7.594819E-5   
1.172758E+3   2.238650E+1   2.238650E+1   2.792660E+1   1.900000E+1   1.900000E+1   0.000000E+0   1.900000E+1   1.900000E+1   5.907784E-2   6.925056E-5   
1.178564E+3   2.239099E+1   2.239099E+1   2.809121E+1   9.000000E+0   9.000000E+0   0.000000E+0   9.000000E+0   9.000000E+0   6.515942E-2   7.471051E-5   
1.184248E+3   2.239391E+1   2.239391E+1   2.792169E+1   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   0.000000E+0   6.602823E-2   7.502197E-5   
1.190074E+3   2.239001E+1   2.239001E+1   2.778790E+1   -9.000000E+0   -9.000000E+0   0.000000E+0   -9.000000E+0   -9.000000E+0   6.255298E-2   7.099136E-5   
1.195980E+3   2.238070E+1   2.238070E+1   2.794430E+1   -1.900000E+1   -1.900000E+1   0.000000E+0   -1.900000E+1   -1.900000E+1   5.994656E-2   6.776730E-5   
1.201915E+3   2.239059E+1   2.239059E+1   2.803411E+1   -2.900000E+1   -2.900000E+1   0.000000E+0   -2.800000E+1   -2.800000E+1   6.689705E-2   7.415765E-5   
1.207799E+3   2.239370E+1   2.239370E+1   2.805041E+1   -3.900000E+1   -3.900000E+1   0.000000E+0   -3.900000E+1   -3.900000E+1   6.602825E-2   7.260853E-5   
1.213706E+3   2.240301E+1   2.240301E+1   2.791021E+1   -4.900000E+1   -4.900000E+1   0.000000E+0   -4.900000E+1   -4.900000E+1   6.602819E-2   7.198964E-5   
1.219637E+3   2.239459E+1   2.239459E+1   2.777169E+1   -5.900000E+1   -5.900000E+1   0.000000E+0   -5.900000E+1   -5.900000E+1   -2.171980E-2   -1.633693E-5   
1.225499E+3   2.240740E+1   2.240740E+1   2.766180E+1   -6.900000E+1   -6.900000E+1   0.000000E+0   -6.900000E+1   -6.900000E+1   -7.645370E-2   -7.166455E-5   
1.231380E+3   2.239871E+1   2.239871E+1   2.765710E+1   -7.900000E+1   -7.900000E+1   0.000000E+0   -7.800000E+1   -7.800000E+1   -9.035434E-2   -8.611576E-5   
1.237258E+3   2.240521E+1   2.240521E+1   2.764211E+1   -8.900000E+1   -8.900000E+1   0.000000E+0   -8.900000E+1   -8.900000E+1   -9.296072E-2   -8.940166E-5   
1.243258E+3   2.240841E+1   2.240841E+1   2.769540E+1   -9.900000E+1   -9.900000E+1   0.000000E+0   -9.900000E+1   -9.900000E+1   -7.906004E-2   -7.612620E-5   
1.260626E+3   2.240820E+1   2.240820E+1   2.766009E+1   -1.500000E+2   -1.500000E+2   0.000000E+0   -1.520000E+2   -1.520000E+2   -8.687918E-2   -8.722158E-5   
1.267805E+3   2.241830E+1   2.241830E+1   2.763021E+1   -1.990000E+2   -1.990000E+2   0.000000E+0   -1.980000E+2   -1.980000E+2   -9.122313E-2   -9.441019E-5   
1.274984E+3   2.242031E+1   2.242031E+1   2.740811E+1   -2.490000E+2   -2.490000E+2   0.000000E+0   -2.480000E+2   -2.480000E+2   -7.645370E-2   -8.274172E-5   
1.282363E+3   2.241299E+1   2.241299E+1   2.735729E+1   -2.990000E+2   -2.990000E+2   0.000000E+0   -2.980000E+2   -2.980000E+2   -8.253523E-2   -9.191464E-5   
1.289553E+3   2.241519E+1   2.241519E+1   2.734680E+1   -3.490000E+2   -3.490000E+2   0.000000E+0   -3.480000E+2   -3.480000E+2   -7.558490E-2   -8.806169E-5   
1.296725E+3   2.241549E+1   2.241549E+1   2.756149E+1   -3.990000E+2   -3.990000E+2   0.000000E+0   -3.980000E+2   -3.980000E+2   -7.819133E-2   -9.376110E-5   
1.303930E+3   2.242239E+1   2.242239E+1   2.749911E+1   -4.490000E+2   -4.490000E+2   0.000000E+0   -4.480000E+2   -4.480000E+2   -7.124093E-2   -8.990808E-5   
1.311077E+3   2.242300E+1   2.242300E+1   2.750939E+1   -4.990000E+2   -4.990000E+2   0.000000E+0   -4.980000E+2   -4.980000E+2   -7.297859E-2   -9.473912E-5   
1.331375E+3   2.241619E+1   2.241619E+1   2.773651E+1   -6.000000E+2   -6.000000E+2   0.000000E+0   -6.020000E+2   -6.020000E+2   -6.689701E-2   -9.509623E-5   
1.339125E+3   2.241940E+1   2.241940E+1   2.769161E+1   -6.990000E+2   -6.990000E+2   0.000000E+0   -6.980000E+2   -6.980000E+2   -5.038991E-2   -8.453753E-5   
1.346981E+3   2.241119E+1   2.241119E+1   2.773150E+1   -7.990000E+2   -7.990000E+2   0.000000E+0   -7.980000E+2   -7.980000E+2   -5.473381E-2   -9.506781E-5   
1.355016E+3   2.240801E+1   2.240801E+1   2.772579E+1   -8.990000E+2   -8.990000E+2   0.000000E+0   -8.980000E+2   -8.980000E+2   -4.604594E-2   -9.257229E-5   
1.362872E+3   2.241079E+1   2.241079E+1   2.776510E+1   -9.990000E+2   -9.990000E+2   0.000000E+0   -9.980000E+2   -9.980000E+2   -3.648931E-2   -8.920842E-5   
1.377182E+3   2.240551E+1   2.240551E+1   2.776101E+1   -1.998000E+3   -1.998000E+3   0.000000E+0   -1.997000E+3   -1.997000E+3   1.911343E-2   -9.545296E-5   
1.389958E+3   2.241921E+1   2.241921E+1   2.791461E+1   -2.998000E+3   -2.998000E+3   0.000000E+0   -2.998000E+3   -2.998000E+3   9.382951E-2   -8.271672E-5   
1.401760E+3   2.240429E+1   2.240429E+1   2.796569E+1   -3.998000E+3   -3.998000E+3   0.000000E+0   -3.997000E+3   -3.997000E+3   1.589889E-1   -7.940902E-5   
1.413043E+3   2.241589E+1   2.241589E+1   2.764889E+1   -4.999000E+3   -4.999000E+3   0.000000E+0   -4.998000E+3   -4.998000E+3   2.145916E-1   -8.577740E-5   
1.425392E+3   2.240829E+1   2.240829E+1   2.762530E+1   -5.999000E+3   -5.999000E+3   0.000000E+0   -5.998000E+3   -5.998000E+3   2.901769E-1   -7.211043E-5   
1.436327E+3   2.240890E+1   2.240890E+1   2.775491E+1   -6.999000E+3   -6.999000E+3   0.000000E+0   -6.997000E+3   -6.997000E+3   3.640237E-1   -6.011923E-5   
1.448125E+3   2.242739E+1   2.242739E+1   2.773931E+1   -7.998000E+3   -7.998000E+3   0.000000E+0   -7.997000E+3   -7.997000E+3   4.248385E-1   -6.121603E-5   
1.460740E+3   2.243041E+1   2.243041E+1   2.782849E+1   -8.999000E+3   -8.999000E+3   0.000000E+0   -8.998000E+3   -8.998000E+3   5.030297E-1   -4.500627E-5   
1.472591E+3   2.241851E+1   2.241851E+1   2.758560E+1   -9.998000E+3   -9.998000E+3   0.000000E+0   -9.997000E+3   -9.997000E+3   5.568958E-1   -5.298666E-5   
1.484207E+3   2.241619E+1   2.241619E+1   2.757781E+1   -1.099900E+4   -1.099900E+4   0.000000E+0   -1.099800E+4   -1.099800E+4   6.281372E-1   -4.372354E-5   
1.497382E+3   2.240341E+1   2.240341E+1   2.770349E+1   -1.199900E+4   -1.199900E+4   0.000000E+0   -1.199800E+4   -1.199800E+4   6.932958E-1   -4.047845E-5   
1.509476E+3   2.239929E+1   2.239929E+1   2.755139E+1   -1.299900E+4   -1.299900E+4   0.000000E+0   -1.299800E+4   -1.299800E+4   7.654069E-1   -3.028410E-5   
1.522585E+3   2.238830E+1   2.238830E+1   2.770779E+1   -1.399800E+4   -1.399800E+4   0.000000E+0   -1.399700E+4   -1.399700E+4   8.340423E-1   -2.350202E-5   
1.535674E+3   2.237469E+1   2.237469E+1   2.784081E+1   -1.499800E+4   -1.499800E+4   0.000000E+0   -1.499700E+4   -1.499700E+4   9.078841E-1   -1.157773E-5   
1.550305E+3   2.236669E+1   2.236669E+1   2.793401E+1   -1.599800E+4   -1.599800E+4   0.000000E+0   -1.599700E+4   -1.599700E+4   9.634894E-1   -1.747572E-5   
1.565940E+3   2.237780E+1   2.237780E+1   2.763329E+1   -1.699900E+4   -1.699900E+4   0.000000E+0   -1.699800E+4   -1.699800E+4   1.028649E+0   -1.246000E-5   
@@END Data.
@Measurement parameters
                                        Upward Part    Downward part  Average        Parameter 'definition'                  
Hysteresis Loop                                                                      Hysteresis Parameters                   
                                                                                                                             
Hc Oe                                   55.707         -57.150        56.429         Coercive Field: Field at which M//H changes sign
Mr emu                                  -85.196E-6     75.022E-6      80.109E-6      Remanent Magnetization: M at H=0        
S                                       0.805          0.772          0.788          Squareness: Mr/Ms                       
S*                                      0.850          0.809          0.829          1-(Mr/Hc)(1/slope at Hc)                
Ms emu                                  105.840E-6     -97.194E-6     101.517E-6     Saturation Magnetization: maximum M measured
                                                                                                                             

@END Measurement parameters
